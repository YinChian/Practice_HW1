module Clock_Counter(
	input CLK_50,
	input oneHz,
	input reset,
	input testSignal,
	output reg [6:0]
);

	always(posedge CLK_50)
	
endmodule